////////////////////////////////////////////////////////////////////////////////// 
// File Name      : temp.sv
// Project        :
// Encrypt        : NO
// Created On     : 16-12-2022  (DD-MM-YYYY)
// Last Modified  : Friday 16 December 2022 04:12:34 PM IST
// Developers     : eInfochips Ltd.
// Description    : 
// Assumptions    : None
// Limitations    : None
// Known Errors   : None
// Revision       :
//
////////////////////////////////////////////////////////////////////////////////// 
////////////////////////////////////////////////////////////////////////////////// 
//                        Copy right Information
// Copyright (c) 1996-2014 eInfochips Ltd. - All rights reserved.
//
// This file is authored by eInfochips Ltd. and is eInfochips
// Ltd. intellectual property, including the copyrights in all countries
// in the world. This file is provided under a license to use only with all
// other rights, including ownership rights, being retained by eInfochips 
// Ltd.
//
// This file may not be distributed, copied, or reproduced in any manner,
// electronic or otherwise, without the express written consent of
// eInfochips Ltd.
////////////////////////////////////////////////////////////////////////////////// 
//================================================================================


nothing there







////////////////////////////////////////////////////////////////////////////////
// Method name         :
// Parameters passed   : None 
// Returned parameters : None
// Description         :
////////////////////////////////////////////////////////////////////////////////






//---------------------------------------------------------------------------------
// End of File
//---------------------------------------------------------------------------------
////////////////////////////////////////////////////////////////////////////////// 
//                        Copy right Information
// Copyright (c) 1996-2014 eInfochips Ltd. - All rights reserved.
//
// This file is authored by eInfochips Ltd. and is eInfochips
// Ltd. intellectual property, including the copyrights in all countries
// in the world. This file is provided under a license to use only with all
// other rights, including ownership rights, being retained by eInfochips 
// Ltd.
//
// This file may not be distributed, copied, or reproduced in any manner,
// electronic or otherwise, without the express written consent of
// eInfochips Ltd.
////////////////////////////////////////////////////////////////////////////////// 
//================================================================================
